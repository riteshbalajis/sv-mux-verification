
class rstgen;
  task rstgen_t();
    #10 rst=0;
  endtask
endclass